`ifndef DEFINES

`define DEFINES

`define ZF 4
`define CF 5
`define OF 6
`define SF 7

`define DELAY 1

`endif
