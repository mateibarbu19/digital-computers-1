module example(
    output out,
    input in
);

    not(out, in);
	
endmodule
