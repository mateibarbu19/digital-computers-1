module module01(
  output out,
  input in
  );

  not(out, in);

endmodule