/* Constants */
`define BTN_PRESS_THLD         5'b01000
`define BTN_RELEASE_THLD			5'b10110
`define BTN_PRESSED_CYCLES		6'b100000
`define CLK_PERIOD					3
`define TIME_TO_OUTPUT			20
`define SECOND						40