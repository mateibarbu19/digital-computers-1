// Copyright 2018 Darius Neatu <neatudarius@gmail.com>

`include "defines.vh"

module test_alu ();

    /* verilator lint_off UNUSED */
	function tester;
		input        [1024 * 8 - 1 : 0] opname;
		input        [4:0]              opcode;
		input signed [7:0]              expected;
		input signed [7:0]              out;
		input signed [3:0]              A;
		input signed [3:0]              B;

		begin
			if (out == expected) begin
				tester = 1'b1;
				$display("%s(%2d, %2d): OK (out = (%4b%4b))", opname, A, B, out[7:4], out[3:0]);
			end else begin
				tester = 1'bx;
				$display("%s(%2d, %2d): FAILED => (%4b%4b) vs (%4b%4b)", opname, A, B, expected[7:4], expected[3:0], out[7:4], out[3:0]);
			end
		end
	endfunction
    /* verilator lint_on UNUSED */

	// outputs
	wire [7:0] out     ;
	reg  [7:0] expected;

	// Inputs
	reg [4:0] opcode;
	reg [3:0] A     ;
	reg [3:0] B     ;

	// checker
	reg [7:0] respect;


	reg [1024*8-1:0] opname;

	// Instantiate the Unit Under Test (UUT)
	alu #(.NR_BITS(4)) UUT (
		.out(out   ),
		.sel(opcode),
		.in0(A     ),
		.in1(B     )
	);

	initial begin
		$dumpfile("alu_test.vcd");
		$dumpvars(0, test_alu);

		// Initialize Inputs
		opcode = 0;
		A = 0;
		B = 0;
		respect = 0;

		#10;

		// =======================================================
		// =======================================================
		// TEST NAND: A = 0, B = 0
		#10;
		opname = "NAND";
		opcode = 5'd1;
		A = 4'b0000;
		B = 4'b0000;
		expected = 8'b0000_1111;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST NAND: A = 15, B = 15
		#10;
		opname = "NAND";
		opcode = 5'd1;
		A = 4'b1111;
		B = 4'b1111;
		expected = 8'b0000_0000;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST NAND: A = 6, B = 9
		#10;
		opname = "NAND";
		opcode = 5'd1;
		A = 4'b0110;
		B = 4'b1001;
		expected = 8'b0000_1111;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST XOR: A = 0, B = 0
		#10;
		opname = "XOR";
		opcode = 5'd2;
		A = 4'b0000;
		B = 4'b0000;
		expected = 8'b0000_0000;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST XOR: A = 3, B = 7
		#10;
		opname = "XOR";
		opcode = 5'd2;
		A = 4'b0011;
		B = 4'b0111;
		expected = 8'b0000_0100;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST XOR: A = 10, B = 5
		#10;
		opname = "XOR";
		opcode = 5'd2;
		A = 4'b1010;
		B = 4'b0101;
		expected = 8'b0000_1111;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST ADD: A = 0, B = 0
		#10;
		opname = "ADD";
		opcode = 5'd4;
		A = 4'b0000;
		B = 4'b0000;
		expected = 8'b0000_0000;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// =======================================================
		// TEST ADD: A = 1, B = 5
		#10;
		opname = "ADD";
		opcode = 5'd4;
		A = 4'b0001;
		B = 4'b0101;
		expected = 8'b0000_0110;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// =======================================================
		// TEST ADD: A = 5, B = 1
		#10;
		opname = "ADD";
		opcode = 5'd4;
		A = 4'b0101;
		B = 4'b0001;
		expected = 8'b0000_0110;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// =======================================================
		// TEST ADD: A = 6, B = 9
		#10;
		opname = "ADD";
		opcode = 5'd4;
		A = 4'b0110;
		B = 4'b1001;
		expected = 8'b0000_1111;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST ADD: A = 6, B = 6
		#10;
		opname = "ADD";
		opcode = 5'd4;
		A = 4'b0110;
		B = 4'b0110;
		expected = 8'b0000_1100;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// =======================================================
		// TEST SUB: A = 0, B = 0
		#10;
		opname = "SUB";
		opcode = 5'd8;
		A = 4'b0000;
		B = 4'b0000;
		expected = 8'b0000_0000;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// =======================================================
		// TEST SUB: A = 7, B = 5
		#10;
		opname = "SUB";
		opcode = 5'd8;
		A = 4'b0111;
		B = 4'b0101;
		expected = 8'b0000_0010;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST SUB: A = 5, B = 7
		#10;
		opname = "SUB";
		opcode = 5'd8;
		A = 4'b0101;
		B = 4'b0111;
		expected = 8'b0000_1110;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================


		// =======================================================
		// =======================================================
		// TEST SUB: A = 2, B = -2
		#10;
		opname = "SUB";
		opcode = 5'd8;
		A = 4'b0010;
		B = 4'b1110;
		expected = 8'b0000_0100;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================




		// =======================================================
		// =======================================================
		// TEST SUB: A = -2, B = -1
		#10;
		opname = "SUB";
		opcode = 5'd8;
		A = 4'b1110;
		B = 4'b1111;
		expected = 8'b0000_1111;
		#10;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// =======================================================
		// TEST MUL: A = 2, B = 0
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b0010;
		B =      4'b0000;
		expected = 8'b0000_0000;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// TEST MUL: A = 2, B = 1
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b0010;
		B =      4'b0001;
		expected = 8'b0000_0010;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// TEST MUL: A = 2, B = -1
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b0010;
		B =      4'b1111;
		expected = 8'b1111_1110;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// TEST MUL: A = 4, B = 4
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b0100;
		B =      4'b0100;
		expected = 8'b0001_0000;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// TEST MUL: A = 4, B = -4
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b0100;
		B =      4'b1100;
		expected = 8'b1111_0000;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// TEST MUL: A = -4, B = 4
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b1100;
		B =      4'b0100;
		expected = 8'b1111_0000;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================



		// =======================================================
		// TEST MUL: A = -4, B = -4
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b1100;
		B =      4'b1100;
		expected = 8'b0001_0000;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================

		// =======================================================
		// TEST MUL: A = -1, B = -6
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b1111;
		B =      4'b1010;
		expected = 8'b0000_0110;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================

		// =======================================================
		// TEST MUL: A = -1, B = 5
		#10;
		opname = "MUL";
		opcode = 5'd16;
		A =      4'b1111;
		B =      4'b0101;
		expected = 8'b1111_1011;
		#20;
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================

		$display("ALU tests = %2d/25", respect);

		$finish();
	end

endmodule
