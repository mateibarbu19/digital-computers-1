`ifndef STATE_MACHINE

`define STATE_MACHINE

`define STATE_RESET		3'h0
`define STATE_IF		3'h1
`define STATE_ID		3'h2
`define STATE_EX		3'h3
`define STATE_MEM		3'h4
`define STATE_WB		3'h5

`endif
