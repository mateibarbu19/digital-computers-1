module module02(
  output out,
  input in
  );

  assign out = ~in;

endmodule
